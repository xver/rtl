interface top_part0_if ;



endinterface
